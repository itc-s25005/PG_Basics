トップガン,卒業白書,マイノリティ・リポート
タイタニック,レヴェナント,インセプション
トレーニングデイ,マイ・ボディガード,フライト
